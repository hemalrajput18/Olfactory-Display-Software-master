** Profile: "SCHEMATIC1-sim_1"  [ C:\Users\hemal\Documents\GitHub\Olfactory-Display-Software\Circuit Diagrams for Tests\ORCAD\m165d25-PSpiceFiles\SCHEMATIC1\sim_1.sim ] 

** Creating circuit file "sim_1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\hemal\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 400us 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
